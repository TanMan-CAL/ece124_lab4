-- Members: Naman Biyani and Tanmay Shah
-- LS206_T20_LAB4

library ieee;
use ieee.std_logic_1164.all;


entity synchronizer is port (

			clk			: in std_logic;
			reset		: in std_logic;
			din			: in std_logic;
			dout		: out std_logic
  );
 end synchronizer;
 
 
architecture circuit of synchronizer is

	Signal sreg				: std_logic_vector(1 downto 0);

BEGIN

	process(clk)
	begin
		if(rising_edge(clk)) then
			if(reset = '1') then
				sreg(0) <= '0';
				sreg(1) <= '0';
				dout <= sreg(1);
			else
				sreg(0) <= din;
				sreg(1) <= sreg(0);
				dout <= sreg(1);
			end if;
		end if;
	end process;
end;
